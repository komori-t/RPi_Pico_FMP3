/*
 *  TOPPERS/ASP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Advanced Standard Profile Kernel
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: tSIOPortTarget.cdl 1363 2020-01-18 02:16:21Z ertl-komori $
 */

/*
 * シリアルインタフェースドライバのターゲット依存部
 * のコンポーネント記述
 */

/*
 * ボードに関する定義
 */
import_C("RP2040.h");

/*
 * USART用 簡易SIOドライバ
 */
import("tUsart.cdl");

/*
 * シリアルインタフェースドライバのターゲット依存部の本体（シリアルイ
 * ンタフェースドライバとSIOドライバを接続する部分）のセルタイプ
 */
celltype tSIOPortTargetMain {
    /*
     *  シリアルインタフェースドライバとの結合
     */
    [inline]   entry    sSIOPort    eSIOPort;
    [optional] call     siSIOCBR    ciSIOCBR;

    /*
     *  SIOドライバとの結合
     */
    call              sSIOPort    cSIOPort;
    [inline] entry    siSIOCBR    eiSIOCBR;

    /*
     *  割込み要求ライン操作のための結合
     */
    call    sInterruptRequest    cInterruptRequest;
};

/*
 * シリアルインタフェースドライバのターゲット依存部（複合コンポーネン
 * ト）のセルタイプ
 */
[active]
composite tSIOPortTarget {
    /*
     * シリアルインタフェースドライバとの結合
     */
    entry              sSIOPort    eSIOPort;
    [optional] call    siSIOCBR    ciSIOCBR;

    /*
     * 属性の定義
     */
    attr {
        uint32_t base;                   /* ベースアドレス */
        uint32_t index;                  /* USARTインデックス */
        INTNO    interruptNumber;        /* 割込み番号 */
        PRI      isrPriority = 1;        /* ISR優先度 */
        PRI      interruptPriority = -2; /* 割込み優先度 */
    };

    /*
     * SIOドライバ
     */
    cell tUsart Usart {
        base     = composite.base;
        index    = composite.index;
        ciSIOCBR = SIOPortMain.eiSIOCBR;
    };

    /*
     * シリアルインタフェースドライバのターゲット依存部の本体
     */
    cell tSIOPortTargetMain SIOPortMain {
        ciSIOCBR          => composite.ciSIOCBR;
        cSIOPort          = Usart.eSIOPort;
        cInterruptRequest = InterruptRequest.eInterruptRequest;
    };
    composite.eSIOPort => SIOPortMain.eSIOPort;

    /*
     * SIOの割込みサービスルーチンと割込み要求ライン
     */
    cell tISR ISRInstance {
        interruptNumber = composite.interruptNumber;
        isrPriority     = composite.isrPriority;
        ciISRBody       = Usart.eiISR;
    };
    cell tInterruptRequest InterruptRequest {
        interruptNumber   = composite.interruptNumber;
        interruptPriority = composite.interruptPriority;
    };
};

/*
 * シリアルインタフェースドライバのターゲット依存部のプロトタイプ
 */
[prototype]
cell tSIOPortTarget SIOPortTarget1 {
    base            = C_EXP("RP2040_UART0_BASE");
    index           = C_EXP("0");
    interruptNumber = C_EXP("RP2040_UART0_IRQn + 16");
};

[prototype]
cell tSIOPortTarget SIOPortTarget2 {
    base            = C_EXP("RP2040_UART1_BASE");
    index           = C_EXP("1");
    interruptNumber = C_EXP("RP2040_UART1_IRQn + 16");
};
